module zero256(z);
output [255:0] z;
 
assign z = 0; 

endmodule
