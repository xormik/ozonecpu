//------------------------------------------------------------------
//-- Verilog Model for RAM
//--	a Single Port 256 line word RAM w/ Synch Read, Synch Write, Synch Reset
//--		Initializes memory to contents in the file "memory.contents"
//--		where each line in the file represents a line in memory in hexidecimal
//--
//-- 	by Ben Liao
//--	Spring 2003 Computer Science 152
//--
//--	256 word lines (32-bit = word)
//--
//--	in order of precedence of signals:
//--		en, rst, we
//--		which means if en == 0 and rst == 1, nothing happens
//-------------------------------------------------------------------
//timing delay is 1ns, accuracy is 1ps
`timescale 1ns / 1ps

module data_source(addr,clk,di,en,rst,we,do);


//-------------Input Signals---------------------------
input [10:0] addr;
input [31:0] 	di;
input 	clk;
input		en;
input		rst;
input		we;

//-------------Parameter Declarations------------------

parameter	ramDelay = 18;
parameter	RAM_depth = 2048;
parameter 	addr_width = 11;
parameter	RAM_width = 32;

//-------------Output Signals--------------------------
output [31:0]   do;

//-------------Port Declarations-----------------------
wire [addr_width-1:0] 	addr;
wire [RAM_width-1:0] 	di;
wire 	 	clk;
wire		en;
wire		rst;
wire		we;
wire	write0, write1, write2, write3, write4, write5, write6, write7;

wire [RAM_width-1:0]	do;
wire [RAM_width-1:0]	do0;
wire [RAM_width-1:0]	do1;
wire [RAM_width-1:0]	do2;
wire [RAM_width-1:0]	do3;
wire [RAM_width-1:0]	do4;
wire [RAM_width-1:0]	do5;
wire [RAM_width-1:0]	do6;
wire [RAM_width-1:0]	do7;
reg [31:0]	memoryLines 	[0:31];
reg[10:0] addr_reg;
reg tempcount;
//-------------Internal Blocks-------------------------



/***********************************************INITIALIZATION OF RAM***************************************************/


RAMB4_S16 memBlock0h(.WE(write0),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do0[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000240c0c00240d8c1200000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 24c724a6248524642443240225ad258c10208fe1afe025ad258c10288fe13408,INIT_03 = 10248fe125ad258c10238fe125ad258c10228fe1afe7afe6afe5afe4afe3afe2,INIT_04 = 8fe18fe125ad258c10278fe125ad258c10268fe125ad258c10258fe125ad258c,INIT_05 = 258c10258fe125ad258c10248fe125ad258c10238fe125ad258c10228fe10000,INIT_06 = 10228fe1afe1afe18fe18fe18fe125ad258c10278fe125ad258c10268fe125ad,INIT_07 = 8fe18fe18fe1afe5afe6afe725ad258c10248fe125ad258c10238fe125ad258c,INIT_08 = afe1afe1afe4afe3afe225ad258c10258fe125ad258c10268fe125ad258c1027,INIT_09 = afe4afe3afe28fe125ad258c10248fe125ad258c10238fe125ad258c10228fe1,INIT_0A = ac12ac1202728c1325ad258c10258fe125ad258c10258fe1afe1afe7afe6afe5,INIT_0B = 0000000000000000000000000000000000000000000008000000ac0cac0d0000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock0h.INIT_00 =
		256'h0000000000000000000000000000000000000000240c0c00240d8c1200000000;
      defparam memBlock0h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0h.INIT_02 =
      256'h24c724a6248524642443240225ad258c10208fe1afe025ad258c10288fe13408;
      defparam memBlock0h.INIT_03 =
      256'h10248fe125ad258c10238fe125ad258c10228fe1afe7afe6afe5afe4afe3afe2;
      defparam memBlock0h.INIT_04 =
      256'h8fe18fe125ad258c10278fe125ad258c10268fe125ad258c10258fe125ad258c;
      defparam memBlock0h.INIT_05 =
      256'h258c10258fe125ad258c10248fe125ad258c10238fe125ad258c10228fe10000;
      defparam memBlock0h.INIT_06 =
      256'h10228fe1afe1afe18fe18fe18fe125ad258c10278fe125ad258c10268fe125ad;
      defparam memBlock0h.INIT_07 =
      256'h8fe18fe18fe1afe5afe6afe725ad258c10248fe125ad258c10238fe125ad258c;
      defparam memBlock0h.INIT_08 =
      256'hafe1afe1afe4afe3afe225ad258c10258fe125ad258c10268fe125ad258c1027;
      defparam memBlock0h.INIT_09 =
      256'hafe4afe3afe28fe125ad258c10248fe125ad258c10238fe125ad258c10228fe1;
      defparam memBlock0h.INIT_0A =
      256'hac12ac1202728c1325ad258c10258fe125ad258c10258fe1afe1afe7afe6afe5;
      defparam memBlock0h.INIT_0B =
      256'h0000000000000000000000000000000000000000000008000000ac0cac0d0000;
      defparam memBlock0h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock0l(.WE(write0),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do0[15:0]))/* synthesis  
xc_props="INIT_00 = 000900080007000600050004000300020001f00d0000001e0000fffc000000b3,INIT_01 = 0019001800170016001500140013001200110010000f000e000d000c000b000a,INIT_02 = 00010001000100010001beef000200010002000000000001000100020000f00d,INIT_03 = 0002000c00040001000200080004000100020004001800140010000c00080004,INIT_04 = 2020200000040001000200180004000100020014000400010002001000040001,INIT_05 = 000100020010000800010002000c0008000100020008000800010002000403cd,INIT_06 = 0002000424082000000800040000000800010002001800080001000200140008,INIT_07 = 200000200000200820042000001000010002000c001000010002000800100001,INIT_08 = 0020000020082004200000200001000220080020000100022004002000010002,INIT_09 = 2004200420042004004000010002200800400001000220040040000100022000,INIT_0A = fff0fff49023fffc008000010002200400800001000220042000200020002004,INIT_0B = 0000000000000000000000000000000000000000000000af024dfff0fff4004d,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock0l.INIT_00 =
		256'h000900080007000600050004000300020001f00d0000001e0000fffc000000b3;
      defparam memBlock0l.INIT_01 =
      256'h0019001800170016001500140013001200110010000f000e000d000c000b000a;
      defparam memBlock0l.INIT_02 =
      256'h00010001000100010001beef000200010002000000000001000100020000f00d;
      defparam memBlock0l.INIT_03 =
      256'h0002000c00040001000200080004000100020004001800140010000c00080004;
      defparam memBlock0l.INIT_04 =
      256'h2020200000040001000200180004000100020014000400010002001000040001;
      defparam memBlock0l.INIT_05 =
      256'h000100020010000800010002000c0008000100020008000800010002000403cd;
      defparam memBlock0l.INIT_06 =
      256'h0002000424082000000800040000000800010002001800080001000200140008;
      defparam memBlock0l.INIT_07 =
      256'h200000200000200820042000001000010002000c001000010002000800100001;
      defparam memBlock0l.INIT_08 =
      256'h0020000020082004200000200001000220080020000100022004002000010002;
      defparam memBlock0l.INIT_09 =
      256'h2004200420042004004000010002200800400001000220040040000100022000;
      defparam memBlock0l.INIT_0A =
      256'hfff0fff49023fffc008000010002200400800001000220042000200020002004;
      defparam memBlock0l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000af024dfff0fff4004d;
      defparam memBlock0l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock0l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock1h(.WE(write1),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do1[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock1h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock1l(.WE(write1),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do1[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock1l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock1l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock2h(.WE(write2),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do2[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock2h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock2l(.WE(write2),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do2[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock2l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock2l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock3h(.WE(write3),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do3[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock3h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock3l(.WE(write3),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do3[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock3l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock3l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock4h(.WE(write4),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do4[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock4h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock4l(.WE(write4),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do4[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock4l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock4l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock5h(.WE(write5),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do5[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock5h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock5l(.WE(write5),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do5[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock5l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock5l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock6h(.WE(write6),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do6[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock6h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock6l(.WE(write6),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do6[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock6l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock6l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock7h(.WE(write7),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[31:16]),.DO(do7[31:16]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock7h.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7h.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on
RAMB4_S16 memBlock7l(.WE(write7),.EN(en),.RST(rst),.CLK(clk),.ADDR(addr[7:0]),.DI(di[15:0]),.DO(do7[15:0]))/* synthesis  
xc_props="INIT_00 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_01 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_02 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_03 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_04 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_05 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_07 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_08 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_09 = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0A = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0B = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0C = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0D = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0E = 0000000000000000000000000000000000000000000000000000000000000000,INIT_0F = 0000000000000000000000000000000000000000000000000000000000000000"*/;
	// synthesis translate_off
		defparam memBlock7l.INIT_00 =
		256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_01 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_02 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_03 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_04 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_05 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_06 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_07 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_08 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_09 =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0A =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0B =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0C =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0D =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0E =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
      defparam memBlock7l.INIT_0F =
      256'h0000000000000000000000000000000000000000000000000000000000000000;
  // synthesis translate_on





//-------------Module Behavior-------------------------
//Initialize Memory contents to the file memory.contents
assign write0 = ((en == 1) && (we == 1)&& (addr[10:8]==0))? 1:0;
assign write1 = ((en == 1) && (we == 1)&& (addr[10:8]==1))? 1:0;
assign write2 = ((en == 1) && (we == 1)&& (addr[10:8]==2))? 1:0;
assign write3 = ((en == 1) && (we == 1)&& (addr[10:8]==3))? 1:0;
assign write4 = ((en == 1) && (we == 1)&& (addr[10:8]==4))? 1:0;
assign write5 = ((en == 1) && (we == 1)&& (addr[10:8]==5))? 1:0;
assign write6 = ((en == 1) && (we == 1)&& (addr[10:8]==6))? 1:0;
assign write7 = ((en == 1) && (we == 1)&& (addr[10:8]==7))? 1:0;

always @(posedge clk) begin
	      addr_reg <= addr;
	   end

assign do = (addr_reg[10:8] == 0)? do0 :
				(addr_reg[10:8] == 1)? do1 :
				(addr_reg[10:8] == 2)? do2 :
(addr_reg[10:8] == 3)? do3 :
				(addr_reg[10:8] == 4)? do4 :
				(addr_reg[10:8] == 5)? do5 :
				(addr_reg[10:8] == 6)? do6 :
				(addr_reg[10:8] == 7)? do7: 0;

endmodule
