module four(four);
	output [31:0] four;

	assign four = 32'd4;
endmodule
