/** Instruction Fetch Unit
 *  Author: Richard Lin
 */

module IFetch();

endmodule
