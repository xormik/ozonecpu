module start_addr(startAddr);

  output [31:0] startAddr;

  assign startAddr = 32'hFFFFFF00;

endmodule




