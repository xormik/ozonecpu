// Arbitrates access to the Common Data Bus
// Basic Operation:  

module CDBArbiter();

  input clk, rst;
  
  // request signals (from each functional unit and buffer)

  // request granted signals (to each functional unit and buffer)

  always @ (posedge clk)
  begin

  // ptr to each request signal?


  end

endmodule
