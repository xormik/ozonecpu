module Zeroes(zeroesO);
output [33:0] zeroesO;
 
assign zeroesO = 34'b0; 

endmodule
