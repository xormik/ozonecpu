module MultDivid_divisor_multiplier_posTwo(in0,out0);
    input [33:0] in0;
    output [33:0] out0;

	 assign out0 = in0  << 1;

endmodule

